package FirstAttempt
    // my first bsv program of the year
endpackage
