`define lambda(arg, body) begin function absolutely_unlikely_name(arg)\
   = body; absolutely_unlikely_name; end
