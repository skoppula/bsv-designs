`define use(pac) import pac::*; export pac::*;

// Standard BSV modules
`use(Assert)
`use(ClientServer)
`use(Clocks)
`use(Connectable)
`use(FIFO)
`use(FIFOF)
`use(FShow)
`use(GetPut)
`use(List)
`use(NumberTypes)
`use(RegFile)
`use(SpecialFIFOs)
`use(StmtFSM)
`use(Vector)

// Extensions
`use(AReg)
`use(AV)
`use(Credit)
`use(Ehr)
`use(GetPutClientServer)
`use(ListOps)
`use(MiscFunctions)
`use(MiscModules)
`use(TAddr)
`use(Trace)
`use(VectorOps)
`use(Abbrevs)
`use(EqCheck)
`use(Loop)

`undef use
